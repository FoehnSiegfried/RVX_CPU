`include "RVX_Info.v"

module Unit_Stage_WD (
    input wire clk,
    input wire rst
);
    
endmodule